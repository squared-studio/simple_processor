/*
Write a markdown documentation for this systemverilog module:
Author : Shahid Uddin Ahmed (shahidshakib0@gmail.com)
*/

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-LOCALPARAMS GENERATED
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-TYPEDEFS
  //////////////////////////////////////////////////////////////////////////////////////////////////
  
  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SIGNALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

`include "sp_pkg.sv"//INCLUDE BECAUSE NO FLIST PRESENT
module instruction_decoder
  import sp_pkg::*;//-PACKAGES//-PARAMETERS //-LOCALPARAMS
(
    input  logic  [          ILEN-1:0] code_i,// INPUT INSTRUCTUIN CODE, ILEN = 16 BIT
    output logic                       func_valid_o,// VALID, 0 OR 1
    output func_t                      func_o,//OPPCODE, ENUM TYPEDEF 
    output logic  [REG_ADDR_WIDTH-1:0] rd_o,//DESTINATION REGISTER, REG_ADD_WIDTH = 3 BIT
    output logic  [REG_ADDR_WIDTH-1:0] rs1_o,// SOURCE REGISTER 1
    output logic  [REG_ADDR_WIDTH-1:0] rs2_o,//SOURCE REGISTER 2
    output logic  [          XLEN-1:0] imm_o//IMMEDIATE VALUE, XLEN = 32 BIT
);
  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-ASSIGNMENTS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  assign rd_o = code_i[15:13];//ADDRESS BIT 13 TO 15 FOR DESTINATION REGISTER
  assign rs1_o = code_i[12:10];//ADDRESS BIT 10 TO 12 FOR SOURCE REGISTER 1
  assign rs2_o = code_i[9:7];//ADDRESS BIT 7 TO 9 FOR SOURCE REGISTER 2
  assign imm_o[5:0] = code_i[9:4];//ADDRESS BIT 4 TO 9 FOR IMMEDIATE VALUE
  assign imm_o[31:6] = code_i[9] ? '1 : '0;//REMAIN 26 BIT WILL BE FILLED WITH THE MSB OF IMMEDIATE VALUE
  
  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-RTLS
  //////////////////////////////////////////////////////////////////////////////////////////////////
  
  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-METHODS
  //////////////////////////////////////////////////////////////////////////////////////////////////
  
  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SEQUENTIALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-INITIAL CHECKS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-COMBINATIONAL
  //////////////////////////////////////////////////////////////////////////////////////////////////

  always_comb begin//COMBINATIONAL BLOCK
    case (code_i[3:0])//CASE WHERE OPCODE 
      default: begin func_o = INVAL; func_valid_o = '0; end//VALID = 0 FOR DEFAULT VALUE OR INVALID VALUE 
      'b0001:  begin func_o = ADDI ; func_valid_o = '1; end//RD = RS1 + IMM
      'b0011:  begin func_o = ADD  ; func_valid_o = '1; end//RD = RS1 + RS2
      'b1011:  begin func_o = SUB  ; func_valid_o = '1; end//RD = RS1 - RS2
      'b0101:  begin func_o = AND  ; func_valid_o = '1; end//RD = RS1 & RS2
      'b1101:  begin func_o = OR   ; func_valid_o = '1; end//RD = RS1 | RS2
      'b1111:  begin func_o = XOR  ; func_valid_o = '1; end//RD = RS1 ^ RS2
      'b0111:  begin func_o = NOT  ; func_valid_o = '1; end//RD = ~RS1
      'b0010:  begin func_o = LOAD ; func_valid_o = '1; end//RD = mem[RS1]
      'b1010:  begin func_o = STORE; func_valid_o = '1; end//mem[RS1] = RS2
      'b0110:  begin func_o = SLL  ; func_valid_o = '1; end//RD = RS1 >> RS2
      'b0100:  begin func_o = SLR  ; func_valid_o = '1; end//RD = RS1 << RS2
      'b1110:  begin func_o = SLLI ; func_valid_o = '1; end//RD = RS1 >> IMM
      'b1100:  begin func_o = SLRI ; func_valid_o = '1; end//RD = RS1 << IMM
    endcase
  end
  
//   `ifdef SIMULATION
//   initial begin
//     if (DATA_WIDTH > 2) begin
//       $display("\033[1;33m%m DATA_WIDTH\033[0m");
//     end
//   end
// `endif  // SIMULATION

endmodule




  
  
  

  

  

  



